** sch_path: /home/anton/projects/tt-vga-fun/xschem/b.sch
**.subckt b
V1 vramp GND pwl 0ns 0v, 20ns 0v, 100ns 1.8v, 200ns 1.8v
V2 vpwr GND 1.8
V3 v040n GND pulse 1.8v 0v 0n 1n 1n 19n 40n
V4 v080n GND pulse 1.8v 0v 0n 1n 1n 39n 80n
V5 v160n GND pulse 1.8v 0v 0n 1n 1n 79n 160n
x5 vdac4pin vdac4 GND tt06_analog_load
R8 vdac4pin GND 1e6 m=1
V6 v320n GND pulse 1.8v 0v 0n 1n 1n 159n 320n
V7 v640n GND pulse 1.8v 0v 0n 1n 1n 319n 640n
V8 v1280n GND pulse 1.8v 0v 0n 1n 1n 639n 1280n
V9 v2560n GND pulse 1.8v 0v 0n 1n 1n 1279n 2560n
V10 v5120n GND pulse 1.8v 0v 0n 1n 1n 2559n 5120n
x7 vpwr GND v040n v080n v160n v320n v640n v1280n v2560n v5120n vdac4 bdac
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/anton/.volare/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/anton/.volare/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/anton/.volare/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/anton/.volare/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice





.options savecurrents

.control
  save all
  tran 1n 6400n
  write b.raw
*  plot
*  + i(vsteer)
*  plot
*  + vdac1 vdac2 vdac3


  plot
  + vdac4*30 vdac4pin*30
  + v040n+2.0
  + v080n+4
  + v160n+6
  + v320n+8
  + v640n+10
  + v1280n+12
  + v2560n+14
  + v5120n+16
*v5120n/2.0 + v2560n/4.0 + v1280n/8.0 + v640n/16.0 + v320n/32.0 + v160n/64.0 + v080n/128.0 + v040n/256.0


*  plot vpull
*  + vramp
*  + v040n
*  + v080n+2
*  + v160n+4
.endc




**** end user architecture code
**.ends

* expanding   symbol:  tt06_analog_load.sym # of pins=3
** sym_path: /home/anton/projects/tt-vga-fun/xschem/tt06_analog_load.sym
** sch_path: /home/anton/projects/tt-vga-fun/xschem/tt06_analog_load.sch
.subckt tt06_analog_load a_ext a_int GND
*.iopin a_int
*.iopin a_ext
*.iopin GND
R1 a_ext a_int 500 m=1
C1 a_int GND 2.5p m=1
C2 a_ext GND 2.5p m=1
.ends


* expanding   symbol:  bdac.sym # of pins=11
** sym_path: /home/anton/projects/tt-vga-fun/xschem/bdac.sym
** sch_path: /home/anton/projects/tt-vga-fun/xschem/bdac.sch
.subckt bdac vcc vss d0 d1 d2 d3 d4 d5 d6 d7 vdac
*.ipin d0
*.opin vdac
*.iopin vcc
*.ipin d1
*.ipin d2
*.ipin d3
*.ipin d4
*.ipin d5
*.ipin d6
*.ipin d7
*.iopin vss
XM1 net5 net2 net1 net1 sky130_fd_pr__pfet_01v8 L=1 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 net4 net2 net1 net1 sky130_fd_pr__pfet_01v8 L=2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 net3 net2 net1 net1 sky130_fd_pr__pfet_01v8 L=4 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 net2 net2 net1 net1 sky130_fd_pr__pfet_01v8 L=0.5 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net3 d0 vdac vdac sky130_fd_pr__nfet_01v8 L=2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 net4 d1 vdac vdac sky130_fd_pr__nfet_01v8 L=1.2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 net5 d2 vdac vdac sky130_fd_pr__nfet_01v8 L=0.5 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 vdac vcc vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 net6 net2 net1 net1 sky130_fd_pr__pfet_01v8 L=0.5 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 net6 d3 vdac vdac sky130_fd_pr__nfet_01v8 L=0.25 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM11 net7 net2 net1 net1 sky130_fd_pr__pfet_01v8 L=0.25 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM12 net7 d4 vdac vdac sky130_fd_pr__nfet_01v8 L=0.6 W=0.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM13 net8 net2 net1 net1 sky130_fd_pr__pfet_01v8 L=0.3 W=1.35 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM14 net8 d5 vdac vdac sky130_fd_pr__nfet_01v8 L=0.25 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM15 net9 net2 net1 net1 sky130_fd_pr__pfet_01v8 L=0.25 W=2.1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM16 net9 d6 vdac vdac sky130_fd_pr__nfet_01v8 L=0.25 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM17 net10 net2 net1 net1 sky130_fd_pr__pfet_01v8 L=0.25 W=4.3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM18 net10 d7 vdac vdac sky130_fd_pr__nfet_01v8 L=0.15 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM19 net2 vcc vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XR5 net1 vcc vss sky130_fd_pr__res_high_po_5p73 L=10 mult=1 m=1
XM20 net11 vcc vss vss sky130_fd_pr__nfet_01v8 L=0.6 W=10 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XC1 net11 vdac sky130_fd_pr__cap_mim_m3_1 W=28 L=20 MF=1 m=1
.ends

.GLOBAL GND
.end
